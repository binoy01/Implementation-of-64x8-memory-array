magic
tech sky130B
magscale 1 2
timestamp 1658299083
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 3698 119200 3754 120000
rect 5998 119200 6054 120000
rect 8298 119200 8354 120000
rect 10598 119200 10654 120000
rect 12898 119200 12954 120000
rect 15198 119200 15254 120000
rect 17498 119200 17554 120000
rect 19798 119200 19854 120000
rect 22098 119200 22154 120000
rect 24398 119200 24454 120000
rect 26698 119200 26754 120000
rect 28998 119200 29054 120000
rect 31298 119200 31354 120000
rect 33598 119200 33654 120000
rect 35898 119200 35954 120000
rect 38198 119200 38254 120000
rect 40498 119200 40554 120000
rect 42798 119200 42854 120000
rect 45098 119200 45154 120000
rect 47398 119200 47454 120000
rect 49698 119200 49754 120000
rect 51998 119200 52054 120000
rect 54298 119200 54354 120000
rect 56598 119200 56654 120000
rect 58898 119200 58954 120000
rect 61198 119200 61254 120000
rect 63498 119200 63554 120000
rect 65798 119200 65854 120000
rect 68098 119200 68154 120000
rect 70398 119200 70454 120000
rect 72698 119200 72754 120000
rect 74998 119200 75054 120000
rect 77298 119200 77354 120000
rect 79598 119200 79654 120000
rect 81898 119200 81954 120000
rect 84198 119200 84254 120000
rect 86498 119200 86554 120000
rect 88798 119200 88854 120000
rect 91098 119200 91154 120000
rect 93398 119200 93454 120000
rect 95698 119200 95754 120000
rect 97998 119200 98054 120000
rect 100298 119200 100354 120000
rect 102598 119200 102654 120000
rect 104898 119200 104954 120000
rect 107198 119200 107254 120000
rect 109498 119200 109554 120000
rect 111798 119200 111854 120000
rect 114098 119200 114154 120000
rect 116398 119200 116454 120000
rect 118698 119200 118754 120000
rect 120998 119200 121054 120000
rect 123298 119200 123354 120000
rect 125598 119200 125654 120000
rect 127898 119200 127954 120000
rect 130198 119200 130254 120000
rect 132498 119200 132554 120000
rect 134798 119200 134854 120000
rect 137098 119200 137154 120000
rect 139398 119200 139454 120000
rect 141698 119200 141754 120000
rect 143998 119200 144054 120000
rect 146298 119200 146354 120000
rect 148598 119200 148654 120000
rect 150898 119200 150954 120000
rect 153198 119200 153254 120000
rect 155498 119200 155554 120000
rect 157798 119200 157854 120000
rect 160098 119200 160154 120000
rect 162398 119200 162454 120000
rect 164698 119200 164754 120000
rect 166998 119200 167054 120000
rect 169298 119200 169354 120000
rect 171598 119200 171654 120000
rect 173898 119200 173954 120000
rect 176198 119200 176254 120000
rect 3146 0 3202 800
rect 8574 0 8630 800
rect 14002 0 14058 800
rect 19430 0 19486 800
rect 24858 0 24914 800
rect 30286 0 30342 800
rect 35714 0 35770 800
rect 41142 0 41198 800
rect 46570 0 46626 800
rect 51998 0 52054 800
rect 57426 0 57482 800
rect 62854 0 62910 800
rect 68282 0 68338 800
rect 73710 0 73766 800
rect 79138 0 79194 800
rect 84566 0 84622 800
rect 89994 0 90050 800
rect 95422 0 95478 800
rect 100850 0 100906 800
rect 106278 0 106334 800
rect 111706 0 111762 800
rect 117134 0 117190 800
rect 122562 0 122618 800
rect 127990 0 128046 800
rect 133418 0 133474 800
rect 138846 0 138902 800
rect 144274 0 144330 800
rect 149702 0 149758 800
rect 155130 0 155186 800
rect 160558 0 160614 800
rect 165986 0 166042 800
rect 171414 0 171470 800
rect 176842 0 176898 800
<< obsm2 >>
rect 3148 119144 3642 119354
rect 3810 119144 5942 119354
rect 6110 119144 8242 119354
rect 8410 119144 10542 119354
rect 10710 119144 12842 119354
rect 13010 119144 15142 119354
rect 15310 119144 17442 119354
rect 17610 119144 19742 119354
rect 19910 119144 22042 119354
rect 22210 119144 24342 119354
rect 24510 119144 26642 119354
rect 26810 119144 28942 119354
rect 29110 119144 31242 119354
rect 31410 119144 33542 119354
rect 33710 119144 35842 119354
rect 36010 119144 38142 119354
rect 38310 119144 40442 119354
rect 40610 119144 42742 119354
rect 42910 119144 45042 119354
rect 45210 119144 47342 119354
rect 47510 119144 49642 119354
rect 49810 119144 51942 119354
rect 52110 119144 54242 119354
rect 54410 119144 56542 119354
rect 56710 119144 58842 119354
rect 59010 119144 61142 119354
rect 61310 119144 63442 119354
rect 63610 119144 65742 119354
rect 65910 119144 68042 119354
rect 68210 119144 70342 119354
rect 70510 119144 72642 119354
rect 72810 119144 74942 119354
rect 75110 119144 77242 119354
rect 77410 119144 79542 119354
rect 79710 119144 81842 119354
rect 82010 119144 84142 119354
rect 84310 119144 86442 119354
rect 86610 119144 88742 119354
rect 88910 119144 91042 119354
rect 91210 119144 93342 119354
rect 93510 119144 95642 119354
rect 95810 119144 97942 119354
rect 98110 119144 100242 119354
rect 100410 119144 102542 119354
rect 102710 119144 104842 119354
rect 105010 119144 107142 119354
rect 107310 119144 109442 119354
rect 109610 119144 111742 119354
rect 111910 119144 114042 119354
rect 114210 119144 116342 119354
rect 116510 119144 118642 119354
rect 118810 119144 120942 119354
rect 121110 119144 123242 119354
rect 123410 119144 125542 119354
rect 125710 119144 127842 119354
rect 128010 119144 130142 119354
rect 130310 119144 132442 119354
rect 132610 119144 134742 119354
rect 134910 119144 137042 119354
rect 137210 119144 139342 119354
rect 139510 119144 141642 119354
rect 141810 119144 143942 119354
rect 144110 119144 146242 119354
rect 146410 119144 148542 119354
rect 148710 119144 150842 119354
rect 151010 119144 153142 119354
rect 153310 119144 155442 119354
rect 155610 119144 157742 119354
rect 157910 119144 160042 119354
rect 160210 119144 162342 119354
rect 162510 119144 164642 119354
rect 164810 119144 166942 119354
rect 167110 119144 169242 119354
rect 169410 119144 171542 119354
rect 171710 119144 173842 119354
rect 174010 119144 176142 119354
rect 176310 119144 176896 119354
rect 3148 856 176896 119144
rect 3258 800 8518 856
rect 8686 800 13946 856
rect 14114 800 19374 856
rect 19542 800 24802 856
rect 24970 800 30230 856
rect 30398 800 35658 856
rect 35826 800 41086 856
rect 41254 800 46514 856
rect 46682 800 51942 856
rect 52110 800 57370 856
rect 57538 800 62798 856
rect 62966 800 68226 856
rect 68394 800 73654 856
rect 73822 800 79082 856
rect 79250 800 84510 856
rect 84678 800 89938 856
rect 90106 800 95366 856
rect 95534 800 100794 856
rect 100962 800 106222 856
rect 106390 800 111650 856
rect 111818 800 117078 856
rect 117246 800 122506 856
rect 122674 800 127934 856
rect 128102 800 133362 856
rect 133530 800 138790 856
rect 138958 800 144218 856
rect 144386 800 149646 856
rect 149814 800 155074 856
rect 155242 800 160502 856
rect 160670 800 165930 856
rect 166098 800 171358 856
rect 171526 800 176786 856
<< obsm3 >>
rect 4210 2143 173486 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal2 s 3698 119200 3754 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 49698 119200 49754 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 54298 119200 54354 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 58898 119200 58954 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 63498 119200 63554 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 68098 119200 68154 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 72698 119200 72754 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 77298 119200 77354 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 81898 119200 81954 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 86498 119200 86554 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 91098 119200 91154 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8298 119200 8354 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 95698 119200 95754 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 100298 119200 100354 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104898 119200 104954 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 109498 119200 109554 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 114098 119200 114154 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 118698 119200 118754 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 123298 119200 123354 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 127898 119200 127954 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 132498 119200 132554 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 137098 119200 137154 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 12898 119200 12954 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 141698 119200 141754 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 146298 119200 146354 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 150898 119200 150954 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 155498 119200 155554 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 160098 119200 160154 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 164698 119200 164754 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 169298 119200 169354 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 173898 119200 173954 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 17498 119200 17554 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 22098 119200 22154 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 26698 119200 26754 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 31298 119200 31354 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 35898 119200 35954 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 40498 119200 40554 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 45098 119200 45154 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5998 119200 6054 120000 6 io_out[0]
port 39 nsew signal output
rlabel metal2 s 51998 119200 52054 120000 6 io_out[10]
port 40 nsew signal output
rlabel metal2 s 56598 119200 56654 120000 6 io_out[11]
port 41 nsew signal output
rlabel metal2 s 61198 119200 61254 120000 6 io_out[12]
port 42 nsew signal output
rlabel metal2 s 65798 119200 65854 120000 6 io_out[13]
port 43 nsew signal output
rlabel metal2 s 70398 119200 70454 120000 6 io_out[14]
port 44 nsew signal output
rlabel metal2 s 74998 119200 75054 120000 6 io_out[15]
port 45 nsew signal output
rlabel metal2 s 79598 119200 79654 120000 6 io_out[16]
port 46 nsew signal output
rlabel metal2 s 84198 119200 84254 120000 6 io_out[17]
port 47 nsew signal output
rlabel metal2 s 88798 119200 88854 120000 6 io_out[18]
port 48 nsew signal output
rlabel metal2 s 93398 119200 93454 120000 6 io_out[19]
port 49 nsew signal output
rlabel metal2 s 10598 119200 10654 120000 6 io_out[1]
port 50 nsew signal output
rlabel metal2 s 97998 119200 98054 120000 6 io_out[20]
port 51 nsew signal output
rlabel metal2 s 102598 119200 102654 120000 6 io_out[21]
port 52 nsew signal output
rlabel metal2 s 107198 119200 107254 120000 6 io_out[22]
port 53 nsew signal output
rlabel metal2 s 111798 119200 111854 120000 6 io_out[23]
port 54 nsew signal output
rlabel metal2 s 116398 119200 116454 120000 6 io_out[24]
port 55 nsew signal output
rlabel metal2 s 120998 119200 121054 120000 6 io_out[25]
port 56 nsew signal output
rlabel metal2 s 125598 119200 125654 120000 6 io_out[26]
port 57 nsew signal output
rlabel metal2 s 130198 119200 130254 120000 6 io_out[27]
port 58 nsew signal output
rlabel metal2 s 134798 119200 134854 120000 6 io_out[28]
port 59 nsew signal output
rlabel metal2 s 139398 119200 139454 120000 6 io_out[29]
port 60 nsew signal output
rlabel metal2 s 15198 119200 15254 120000 6 io_out[2]
port 61 nsew signal output
rlabel metal2 s 143998 119200 144054 120000 6 io_out[30]
port 62 nsew signal output
rlabel metal2 s 148598 119200 148654 120000 6 io_out[31]
port 63 nsew signal output
rlabel metal2 s 153198 119200 153254 120000 6 io_out[32]
port 64 nsew signal output
rlabel metal2 s 157798 119200 157854 120000 6 io_out[33]
port 65 nsew signal output
rlabel metal2 s 162398 119200 162454 120000 6 io_out[34]
port 66 nsew signal output
rlabel metal2 s 166998 119200 167054 120000 6 io_out[35]
port 67 nsew signal output
rlabel metal2 s 171598 119200 171654 120000 6 io_out[36]
port 68 nsew signal output
rlabel metal2 s 176198 119200 176254 120000 6 io_out[37]
port 69 nsew signal output
rlabel metal2 s 19798 119200 19854 120000 6 io_out[3]
port 70 nsew signal output
rlabel metal2 s 24398 119200 24454 120000 6 io_out[4]
port 71 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 io_out[5]
port 72 nsew signal output
rlabel metal2 s 33598 119200 33654 120000 6 io_out[6]
port 73 nsew signal output
rlabel metal2 s 38198 119200 38254 120000 6 io_out[7]
port 74 nsew signal output
rlabel metal2 s 42798 119200 42854 120000 6 io_out[8]
port 75 nsew signal output
rlabel metal2 s 47398 119200 47454 120000 6 io_out[9]
port 76 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 78 nsew ground bidirectional
rlabel metal2 s 3146 0 3202 800 6 wb_clk_i
port 79 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[0]
port 80 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_o[10]
port 81 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 wbs_dat_o[11]
port 82 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 wbs_dat_o[12]
port 83 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 wbs_dat_o[13]
port 84 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 wbs_dat_o[14]
port 85 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 wbs_dat_o[15]
port 86 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 wbs_dat_o[16]
port 87 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 wbs_dat_o[17]
port 88 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 wbs_dat_o[18]
port 89 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 wbs_dat_o[19]
port 90 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[1]
port 91 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 wbs_dat_o[20]
port 92 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 wbs_dat_o[21]
port 93 nsew signal output
rlabel metal2 s 127990 0 128046 800 6 wbs_dat_o[22]
port 94 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 wbs_dat_o[23]
port 95 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 wbs_dat_o[24]
port 96 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 wbs_dat_o[25]
port 97 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 wbs_dat_o[26]
port 98 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 wbs_dat_o[27]
port 99 nsew signal output
rlabel metal2 s 160558 0 160614 800 6 wbs_dat_o[28]
port 100 nsew signal output
rlabel metal2 s 165986 0 166042 800 6 wbs_dat_o[29]
port 101 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[2]
port 102 nsew signal output
rlabel metal2 s 171414 0 171470 800 6 wbs_dat_o[30]
port 103 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 wbs_dat_o[31]
port 104 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_o[3]
port 105 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[4]
port 106 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[5]
port 107 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[6]
port 108 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_o[7]
port 109 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 wbs_dat_o[8]
port 110 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 wbs_dat_o[9]
port 111 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6734454
string GDS_FILE /media/bn/0FDFA1F87CD9FC5A/Implementation-of-8x64-memory-array/openlane/simple/runs/22_07_20_12_04/results/signoff/simple.magic.gds
string GDS_START 315570
<< end >>

